`timescale 1ns / 1ps

module tb_singleRAM();

    reg i_clk;
    reg i_ce;
    reg i_we;
    reg [5:0] i_addr;
    reg [7:0] i_data;

    wire [7:0] o_data;

    singleRAM dut(
        .i_clk(i_clk),
        .i_ce(i_ce),
        .i_we(i_we),
        .i_addr(i_addr),
        .i_data(i_data),

        .o_data(o_data)
    );

    always #5 i_clk = ~i_clk;

    initial begin
        #00 i_clk = 0; i_ce = 0; i_we = 0; i_addr = 0; i_data = 0;
        #20 i_ce = 1; i_we = 1;

        for (integer i= 0; i < 64; i = i + 1) begin
            #20 i_addr = i; i_data = i + 1;
        end       
        
        
        for (integer i = 0; i < 64; i = i + 1) begin
            #20 i_we = 0; i_addr = i;
        end
        #20 $finish;
    end


endmodule
